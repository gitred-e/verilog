module and_d(
    output y,
    input a,b
);
assign y = a & b;
endmodule
